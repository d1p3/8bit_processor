library verilog;
use verilog.vl_types.all;
entity adder_with_overflow_vlg_vec_tst is
end adder_with_overflow_vlg_vec_tst;
