library verilog;
use verilog.vl_types.all;
entity ControlUnit_vlg_check_tst is
    port(
        c0              : in     vl_logic;
        c2              : in     vl_logic;
        c3              : in     vl_logic;
        c4              : in     vl_logic;
        c7              : in     vl_logic;
        c8              : in     vl_logic;
        c9              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ControlUnit_vlg_check_tst;
