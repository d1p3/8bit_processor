library verilog;
use verilog.vl_types.all;
entity pi_po_register_74175_vlg_vec_tst is
end pi_po_register_74175_vlg_vec_tst;
