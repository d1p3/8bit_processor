library verilog;
use verilog.vl_types.all;
entity FourBitUpCounter_vlg_vec_tst is
end FourBitUpCounter_vlg_vec_tst;
